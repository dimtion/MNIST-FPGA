library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity testbench_Ram_W_3 is 
end entity;

architecture tb_ram_3 of testbench_Ram_W_3 is 

begin


end tb_ram_3;
